class boot_c;

    task body();
        #10000ns;
        $display("[ti] this is boot");
    endtask 

endclass
