DWC_pcie_ctrl_x2_dbi_araddr
DWC_pcie_ctrl_x2_dbi_arburst
DWC_pcie_ctrl_x2_dbi_arcache
DWC_pcie_ctrl_x2_dbi_arid
DWC_pcie_ctrl_x2_dbi_arlen
DWC_pcie_ctrl_x2_dbi_arlock
DWC_pcie_ctrl_x2_dbi_arprot
DWC_pcie_ctrl_x2_dbi_arqos
DWC_pcie_ctrl_x2_dbi_arsize
DWC_pcie_ctrl_x2_dbi_awaddr
DWC_pcie_ctrl_x2_dbi_awburst
DWC_pcie_ctrl_x2_dbi_awcache
DWC_pcie_ctrl_x2_dbi_awid
DWC_pcie_ctrl_x2_dbi_awlen
DWC_pcie_ctrl_x2_dbi_awlock
DWC_pcie_ctrl_x2_dbi_awprot
DWC_pcie_ctrl_x2_dbi_awqos
DWC_pcie_ctrl_x2_dbi_awsize
DWC_pcie_ctrl_x2_dbi_bid
DWC_pcie_ctrl_x2_dbi_bresp
DWC_pcie_ctrl_x2_dbi_cactive
DWC_pcie_ctrl_x2_dbi_csysack
DWC_pcie_ctrl_x2_dbi_csysreq
DWC_pcie_ctrl_x2_dbi_rdata
DWC_pcie_ctrl_x2_dbi_rid
DWC_pcie_ctrl_x2_dbi_rresp
DWC_pcie_ctrl_x2_dbi_wdata
DWC_pcie_ctrl_x2_dbi_wstrb
DWC_pcie_ctrl_x2_mstr_araddr
DWC_pcie_ctrl_x2_mstr_arburst
DWC_pcie_ctrl_x2_mstr_arcache
DWC_pcie_ctrl_x2_mstr_arid
DWC_pcie_ctrl_x2_mstr_arlen
DWC_pcie_ctrl_x2_mstr_arlock
DWC_pcie_ctrl_x2_mstr_arprot
DWC_pcie_ctrl_x2_mstr_arqos
DWC_pcie_ctrl_x2_mstr_arsize
DWC_pcie_ctrl_x2_mstr_awaddr
DWC_pcie_ctrl_x2_mstr_awburst
DWC_pcie_ctrl_x2_mstr_awcache
DWC_pcie_ctrl_x2_mstr_awid
DWC_pcie_ctrl_x2_mstr_awlen
DWC_pcie_ctrl_x2_mstr_awlock
DWC_pcie_ctrl_x2_mstr_awprot
DWC_pcie_ctrl_x2_mstr_awqos
DWC_pcie_ctrl_x2_mstr_awsize
DWC_pcie_ctrl_x2_mstr_bid
DWC_pcie_ctrl_x2_mstr_bready
DWC_pcie_ctrl_x2_mstr_bresp
DWC_pcie_ctrl_x2_mstr_bvalid
DWC_pcie_ctrl_x2_mstr_cactive
DWC_pcie_ctrl_x2_mstr_csysack
DWC_pcie_ctrl_x2_mstr_csysreq
DWC_pcie_ctrl_x2_mstr_rdata
DWC_pcie_ctrl_x2_mstr_rid
DWC_pcie_ctrl_x2_mstr_rlast
DWC_pcie_ctrl_x2_mstr_rready
DWC_pcie_ctrl_x2_mstr_rresp
DWC_pcie_ctrl_x2_mstr_rvalid
DWC_pcie_ctrl_x2_mstr_wdata
DWC_pcie_ctrl_x2_mstr_wlast
DWC_pcie_ctrl_x2_mstr_wstrb
DWC_pcie_ctrl_x2_slv_araddr
DWC_pcie_ctrl_x2_slv_arburst
DWC_pcie_ctrl_x2_slv_arcache
DWC_pcie_ctrl_x2_slv_arid
DWC_pcie_ctrl_x2_slv_arlen
DWC_pcie_ctrl_x2_slv_arlock
DWC_pcie_ctrl_x2_slv_arprot
DWC_pcie_ctrl_x2_slv_arqos
DWC_pcie_ctrl_x2_slv_arsize
DWC_pcie_ctrl_x2_slv_awaddr
DWC_pcie_ctrl_x2_slv_awburst
DWC_pcie_ctrl_x2_slv_awcache
DWC_pcie_ctrl_x2_slv_awid
DWC_pcie_ctrl_x2_slv_awlen
DWC_pcie_ctrl_x2_slv_awlock
DWC_pcie_ctrl_x2_slv_awprot
DWC_pcie_ctrl_x2_slv_awqos
DWC_pcie_ctrl_x2_slv_awsize
DWC_pcie_ctrl_x2_slv_bid
DWC_pcie_ctrl_x2_slv_bresp
DWC_pcie_ctrl_x2_slv_cactive
DWC_pcie_ctrl_x2_slv_csysack
DWC_pcie_ctrl_x2_slv_csysreq
DWC_pcie_ctrl_x2_slv_rdata
DWC_pcie_ctrl_x2_slv_rid
DWC_pcie_ctrl_x2_slv_rresp
DWC_pcie_ctrl_x2_slv_wdata
DWC_pcie_ctrl_x2_slv_wstrb
DWC_pcie_ctrl_x4_dbi_araddr
DWC_pcie_ctrl_x4_dbi_arburst
DWC_pcie_ctrl_x4_dbi_arcache
DWC_pcie_ctrl_x4_dbi_arid
DWC_pcie_ctrl_x4_dbi_arlen
DWC_pcie_ctrl_x4_dbi_arlock
DWC_pcie_ctrl_x4_dbi_arprot
DWC_pcie_ctrl_x4_dbi_arqos
DWC_pcie_ctrl_x4_dbi_arsize
DWC_pcie_ctrl_x4_dbi_awaddr
DWC_pcie_ctrl_x4_dbi_awburst
DWC_pcie_ctrl_x4_dbi_awcache
DWC_pcie_ctrl_x4_dbi_awid
DWC_pcie_ctrl_x4_dbi_awlen
DWC_pcie_ctrl_x4_dbi_awlock
DWC_pcie_ctrl_x4_dbi_awprot
DWC_pcie_ctrl_x4_dbi_awqos
DWC_pcie_ctrl_x4_dbi_awsize
DWC_pcie_ctrl_x4_dbi_bid
DWC_pcie_ctrl_x4_dbi_bresp
DWC_pcie_ctrl_x4_dbi_cactive
DWC_pcie_ctrl_x4_dbi_csysack
DWC_pcie_ctrl_x4_dbi_csysreq
DWC_pcie_ctrl_x4_dbi_rdata
DWC_pcie_ctrl_x4_dbi_rid
DWC_pcie_ctrl_x4_dbi_rresp
DWC_pcie_ctrl_x4_dbi_wdata
DWC_pcie_ctrl_x4_dbi_wstrb
DWC_pcie_ctrl_x4_mstr_araddr
DWC_pcie_ctrl_x4_mstr_arburst
DWC_pcie_ctrl_x4_mstr_arcache
DWC_pcie_ctrl_x4_mstr_arid
DWC_pcie_ctrl_x4_mstr_arlen
DWC_pcie_ctrl_x4_mstr_arlock
DWC_pcie_ctrl_x4_mstr_arprot
DWC_pcie_ctrl_x4_mstr_arqos
DWC_pcie_ctrl_x4_mstr_arsize
DWC_pcie_ctrl_x4_mstr_awaddr
DWC_pcie_ctrl_x4_mstr_awburst
DWC_pcie_ctrl_x4_mstr_awcache
DWC_pcie_ctrl_x4_mstr_awid
DWC_pcie_ctrl_x4_mstr_awlen
DWC_pcie_ctrl_x4_mstr_awlock
DWC_pcie_ctrl_x4_mstr_awprot
DWC_pcie_ctrl_x4_mstr_awqos
DWC_pcie_ctrl_x4_mstr_awsize
DWC_pcie_ctrl_x4_mstr_bid
DWC_pcie_ctrl_x4_mstr_bready
DWC_pcie_ctrl_x4_mstr_bresp
DWC_pcie_ctrl_x4_mstr_bvalid
DWC_pcie_ctrl_x4_mstr_cactive
DWC_pcie_ctrl_x4_mstr_csysack
DWC_pcie_ctrl_x4_mstr_csysreq
DWC_pcie_ctrl_x4_mstr_rdata
DWC_pcie_ctrl_x4_mstr_rid
DWC_pcie_ctrl_x4_mstr_rlast
DWC_pcie_ctrl_x4_mstr_rready
DWC_pcie_ctrl_x4_mstr_rresp
DWC_pcie_ctrl_x4_mstr_rvalid
DWC_pcie_ctrl_x4_mstr_wdata
DWC_pcie_ctrl_x4_mstr_wlast
DWC_pcie_ctrl_x4_mstr_wstrb
DWC_pcie_ctrl_x4_slv_araddr
DWC_pcie_ctrl_x4_slv_arburst
DWC_pcie_ctrl_x4_slv_arcache
DWC_pcie_ctrl_x4_slv_arid
DWC_pcie_ctrl_x4_slv_arlen
DWC_pcie_ctrl_x4_slv_arlock
DWC_pcie_ctrl_x4_slv_arprot
DWC_pcie_ctrl_x4_slv_arqos
DWC_pcie_ctrl_x4_slv_arsize
DWC_pcie_ctrl_x4_slv_awaddr
DWC_pcie_ctrl_x4_slv_awburst
DWC_pcie_ctrl_x4_slv_awcache
DWC_pcie_ctrl_x4_slv_awid
DWC_pcie_ctrl_x4_slv_awlen
DWC_pcie_ctrl_x4_slv_awlock
DWC_pcie_ctrl_x4_slv_awprot
DWC_pcie_ctrl_x4_slv_awqos
DWC_pcie_ctrl_x4_slv_awsize
DWC_pcie_ctrl_x4_slv_bid
DWC_pcie_ctrl_x4_slv_bresp
DWC_pcie_ctrl_x4_slv_cactive
DWC_pcie_ctrl_x4_slv_csysack
DWC_pcie_ctrl_x4_slv_csysreq
DWC_pcie_ctrl_x4_slv_rdata
DWC_pcie_ctrl_x4_slv_rid
DWC_pcie_ctrl_x4_slv_rresp
DWC_pcie_ctrl_x4_slv_wdata
DWC_pcie_ctrl_x4_slv_wstrb
I_TEST_MODE_PCIE_PHY
PCIE_PHY_APB2CR_QACCEPTn
PCIE_PHY_APB2CR_QACTIVE
PCIE_PHY_APB2CR_QDENY
PCIE_PHY_APB2CR_QREQn
PCIE_PHY_APB2CR_TEST_MODE
PCIE_PHY_APB2CR_TEST_RESETn
PCIE_PHY_APB2CR_paddr
PCIE_PHY_APB2CR_pclk_100
PCIE_PHY_APB2CR_pclk_300
PCIE_PHY_APB2CR_penable
PCIE_PHY_APB2CR_prdata
PCIE_PHY_APB2CR_pready
PCIE_PHY_APB2CR_presetn
PCIE_PHY_APB2CR_psel
PCIE_PHY_APB2CR_pslverr
PCIE_PHY_APB2CR_pwdata
PCIE_PHY_APB2CR_pwrite
PCIE_PHY_ext_pclk_req
PCIE_PHY_pcs_scan_mode
PCIE_PHY_pcs_scan_pclk
PCIE_PHY_pcs_scan_pcs_clk
PCIE_PHY_pcs_scan_pma_clk
PCIE_PHY_pcs_scan_rst
PCIE_PHY_pcs_scan_rx_clk_div
PCIE_PHY_pcs_scan_shift
PCIE_PHY_pcs_scan_shift_cg
PCIE_PHY_phy0_bs_acmode
PCIE_PHY_phy0_bs_actest
PCIE_PHY_phy0_bs_cdr
PCIE_PHY_phy0_bs_ce
PCIE_PHY_phy0_bs_rx_init
PCIE_PHY_phy0_bs_sdr
PCIE_PHY_phy0_bs_tdi
PCIE_PHY_phy0_bs_tdo
PCIE_PHY_phy0_bs_udr
PCIE_PHY_phy0_cr_para_sel
PCIE_PHY_phy0_dtb_out
PCIE_PHY_phy0_jtag_tck
PCIE_PHY_phy0_jtag_tdi
PCIE_PHY_phy0_jtag_tdo
PCIE_PHY_phy0_jtag_tdo_en
PCIE_PHY_phy0_jtag_tms
PCIE_PHY_phy0_jtag_trst_n
PCIE_PHY_phy0_scan_cr_clk
PCIE_PHY_phy0_scan_cr_in
PCIE_PHY_phy0_scan_cr_out
PCIE_PHY_phy0_scan_mode
PCIE_PHY_phy0_scan_mplla_div16p5_clk
PCIE_PHY_phy0_scan_mplla_div16p5_in
PCIE_PHY_phy0_scan_mplla_div16p5_out
PCIE_PHY_phy0_scan_mplla_div33_clk
PCIE_PHY_phy0_scan_mplla_div66_clk
PCIE_PHY_phy0_scan_mplla_div_clk
PCIE_PHY_phy0_scan_mplla_div_in
PCIE_PHY_phy0_scan_mplla_div_out
PCIE_PHY_phy0_scan_mplla_dword_clk
PCIE_PHY_phy0_scan_mplla_dword_in
PCIE_PHY_phy0_scan_mplla_dword_out
PCIE_PHY_phy0_scan_mplla_fb_clk
PCIE_PHY_phy0_scan_mplla_fb_in
PCIE_PHY_phy0_scan_mplla_fb_out
PCIE_PHY_phy0_scan_mplla_oword_clk
PCIE_PHY_phy0_scan_mplla_qword_clk
PCIE_PHY_phy0_scan_mplla_ref_clk
PCIE_PHY_phy0_scan_mplla_ref_in
PCIE_PHY_phy0_scan_mplla_ref_out
PCIE_PHY_phy0_scan_mplla_ssc_clk
PCIE_PHY_phy0_scan_mplla_ssc_in
PCIE_PHY_phy0_scan_mplla_ssc_out
PCIE_PHY_phy0_scan_mplla_word_clk
PCIE_PHY_phy0_scan_mplla_word_in
PCIE_PHY_phy0_scan_mplla_word_out
PCIE_PHY_phy0_scan_mpllb_div_clk
PCIE_PHY_phy0_scan_mpllb_div_in
PCIE_PHY_phy0_scan_mpllb_div_out
PCIE_PHY_phy0_scan_mpllb_dword_clk
PCIE_PHY_phy0_scan_mpllb_dword_in
PCIE_PHY_phy0_scan_mpllb_dword_out
PCIE_PHY_phy0_scan_mpllb_fb_clk
PCIE_PHY_phy0_scan_mpllb_fb_in
PCIE_PHY_phy0_scan_mpllb_fb_out
PCIE_PHY_phy0_scan_mpllb_oword_clk
PCIE_PHY_phy0_scan_mpllb_qword_clk
PCIE_PHY_phy0_scan_mpllb_ref_clk
PCIE_PHY_phy0_scan_mpllb_ref_in
PCIE_PHY_phy0_scan_mpllb_ref_out
PCIE_PHY_phy0_scan_mpllb_ssc_clk
PCIE_PHY_phy0_scan_mpllb_ssc_in
PCIE_PHY_phy0_scan_mpllb_ssc_out
PCIE_PHY_phy0_scan_mpllb_word_clk
PCIE_PHY_phy0_scan_mpllb_word_in
PCIE_PHY_phy0_scan_mpllb_word_out
PCIE_PHY_phy0_scan_phy_ref_dig_clk
PCIE_PHY_phy0_scan_phy_ref_dig_in
PCIE_PHY_phy0_scan_phy_ref_dig_out
PCIE_PHY_phy0_scan_ref_clk
PCIE_PHY_phy0_scan_ref_dig_clk
PCIE_PHY_phy0_scan_ref_dig_in
PCIE_PHY_phy0_scan_ref_dig_out
PCIE_PHY_phy0_scan_ref_in
PCIE_PHY_phy0_scan_ref_out
PCIE_PHY_phy0_scan_ref_range_clk
PCIE_PHY_phy0_scan_ref_range_in
PCIE_PHY_phy0_scan_ref_range_out
PCIE_PHY_phy0_scan_set_rst
PCIE_PHY_phy0_scan_shift
PCIE_PHY_phy0_scan_shift_cg
PCIE_PHY_phy0_sram_bypass
PCIE_PHY_phy0_test_flyover_en
PCIE_PHY_phy_lane0_rx2tx_par_lb_en
PCIE_PHY_phy_lane1_rx2tx_par_lb_en
PCIE_PHY_phy_lane2_rx2tx_par_lb_en
PCIE_PHY_phy_lane3_rx2tx_par_lb_en
PCIE_PHY_phy_reset
PCIE_PHY_phy_rx0_flyover_data_m
PCIE_PHY_phy_rx0_flyover_data_p
PCIE_PHY_phy_rx1_flyover_data_m
PCIE_PHY_phy_rx1_flyover_data_p
PCIE_PHY_phy_rx2_flyover_data_m
PCIE_PHY_phy_rx2_flyover_data_p
PCIE_PHY_phy_rx3_flyover_data_m
PCIE_PHY_phy_rx3_flyover_data_p
PCIE_PHY_phy_scan_rx0_adpt_clk
PCIE_PHY_phy_scan_rx0_adpt_in
PCIE_PHY_phy_scan_rx0_adpt_out
PCIE_PHY_phy_scan_rx0_asic_clk
PCIE_PHY_phy_scan_rx0_asic_in
PCIE_PHY_phy_scan_rx0_asic_out
PCIE_PHY_phy_scan_rx0_div16p5_clk
PCIE_PHY_phy_scan_rx0_div16p5_in
PCIE_PHY_phy_scan_rx0_div16p5_out
PCIE_PHY_phy_scan_rx0_dpll_clk
PCIE_PHY_phy_scan_rx0_dpll_in
PCIE_PHY_phy_scan_rx0_dpll_out
PCIE_PHY_phy_scan_rx0_dword_clk
PCIE_PHY_phy_scan_rx0_dword_in
PCIE_PHY_phy_scan_rx0_dword_out
PCIE_PHY_phy_scan_rx0_scope_clk
PCIE_PHY_phy_scan_rx0_scope_in
PCIE_PHY_phy_scan_rx0_scope_out
PCIE_PHY_phy_scan_rx0_stat_clk
PCIE_PHY_phy_scan_rx0_stat_in
PCIE_PHY_phy_scan_rx0_stat_out
PCIE_PHY_phy_scan_rx0_word_clk
PCIE_PHY_phy_scan_rx0_word_in
PCIE_PHY_phy_scan_rx0_word_out
PCIE_PHY_phy_scan_rx1_adpt_clk
PCIE_PHY_phy_scan_rx1_adpt_in
PCIE_PHY_phy_scan_rx1_adpt_out
PCIE_PHY_phy_scan_rx1_asic_clk
PCIE_PHY_phy_scan_rx1_asic_in
PCIE_PHY_phy_scan_rx1_asic_out
PCIE_PHY_phy_scan_rx1_div16p5_clk
PCIE_PHY_phy_scan_rx1_div16p5_in
PCIE_PHY_phy_scan_rx1_div16p5_out
PCIE_PHY_phy_scan_rx1_dpll_clk
PCIE_PHY_phy_scan_rx1_dpll_in
PCIE_PHY_phy_scan_rx1_dpll_out
PCIE_PHY_phy_scan_rx1_dword_clk
PCIE_PHY_phy_scan_rx1_dword_in
PCIE_PHY_phy_scan_rx1_dword_out
PCIE_PHY_phy_scan_rx1_scope_clk
PCIE_PHY_phy_scan_rx1_scope_in
PCIE_PHY_phy_scan_rx1_scope_out
PCIE_PHY_phy_scan_rx1_stat_clk
PCIE_PHY_phy_scan_rx1_stat_in
PCIE_PHY_phy_scan_rx1_stat_out
PCIE_PHY_phy_scan_rx1_word_clk
PCIE_PHY_phy_scan_rx1_word_in
PCIE_PHY_phy_scan_rx1_word_out
PCIE_PHY_phy_scan_rx2_adpt_clk
PCIE_PHY_phy_scan_rx2_adpt_in
PCIE_PHY_phy_scan_rx2_adpt_out
PCIE_PHY_phy_scan_rx2_asic_clk
PCIE_PHY_phy_scan_rx2_asic_in
PCIE_PHY_phy_scan_rx2_asic_out
PCIE_PHY_phy_scan_rx2_div16p5_clk
PCIE_PHY_phy_scan_rx2_div16p5_in
PCIE_PHY_phy_scan_rx2_div16p5_out
PCIE_PHY_phy_scan_rx2_dpll_clk
PCIE_PHY_phy_scan_rx2_dpll_in
PCIE_PHY_phy_scan_rx2_dpll_out
PCIE_PHY_phy_scan_rx2_dword_clk
PCIE_PHY_phy_scan_rx2_dword_in
PCIE_PHY_phy_scan_rx2_dword_out
PCIE_PHY_phy_scan_rx2_scope_clk
PCIE_PHY_phy_scan_rx2_scope_in
PCIE_PHY_phy_scan_rx2_scope_out
PCIE_PHY_phy_scan_rx2_stat_clk
PCIE_PHY_phy_scan_rx2_stat_in
PCIE_PHY_phy_scan_rx2_stat_out
PCIE_PHY_phy_scan_rx2_word_clk
PCIE_PHY_phy_scan_rx2_word_in
PCIE_PHY_phy_scan_rx2_word_out
PCIE_PHY_phy_scan_rx3_adpt_clk
PCIE_PHY_phy_scan_rx3_adpt_in
PCIE_PHY_phy_scan_rx3_adpt_out
PCIE_PHY_phy_scan_rx3_asic_clk
PCIE_PHY_phy_scan_rx3_asic_in
PCIE_PHY_phy_scan_rx3_asic_out
PCIE_PHY_phy_scan_rx3_div16p5_clk
PCIE_PHY_phy_scan_rx3_div16p5_in
PCIE_PHY_phy_scan_rx3_div16p5_out
PCIE_PHY_phy_scan_rx3_dpll_clk
PCIE_PHY_phy_scan_rx3_dpll_in
PCIE_PHY_phy_scan_rx3_dpll_out
PCIE_PHY_phy_scan_rx3_dword_clk
PCIE_PHY_phy_scan_rx3_dword_in
PCIE_PHY_phy_scan_rx3_dword_out
PCIE_PHY_phy_scan_rx3_scope_clk
PCIE_PHY_phy_scan_rx3_scope_in
PCIE_PHY_phy_scan_rx3_scope_out
PCIE_PHY_phy_scan_rx3_stat_clk
PCIE_PHY_phy_scan_rx3_stat_in
PCIE_PHY_phy_scan_rx3_stat_out
PCIE_PHY_phy_scan_rx3_word_clk
PCIE_PHY_phy_scan_rx3_word_in
PCIE_PHY_phy_scan_rx3_word_out
PCIE_PHY_phy_scan_tx0_ana_dword_clk
PCIE_PHY_phy_scan_tx0_ana_dword_in
PCIE_PHY_phy_scan_tx0_ana_dword_out
PCIE_PHY_phy_scan_tx0_ana_word_clk
PCIE_PHY_phy_scan_tx0_ana_word_in
PCIE_PHY_phy_scan_tx0_ana_word_out
PCIE_PHY_phy_scan_tx0_in
PCIE_PHY_phy_scan_tx0_out
PCIE_PHY_phy_scan_tx1_ana_dword_clk
PCIE_PHY_phy_scan_tx1_ana_dword_in
PCIE_PHY_phy_scan_tx1_ana_dword_out
PCIE_PHY_phy_scan_tx1_ana_word_clk
PCIE_PHY_phy_scan_tx1_ana_word_in
PCIE_PHY_phy_scan_tx1_ana_word_out
PCIE_PHY_phy_scan_tx1_in
PCIE_PHY_phy_scan_tx1_out
PCIE_PHY_phy_scan_tx2_ana_dword_clk
PCIE_PHY_phy_scan_tx2_ana_dword_in
PCIE_PHY_phy_scan_tx2_ana_dword_out
PCIE_PHY_phy_scan_tx2_ana_word_clk
PCIE_PHY_phy_scan_tx2_ana_word_in
PCIE_PHY_phy_scan_tx2_ana_word_out
PCIE_PHY_phy_scan_tx2_in
PCIE_PHY_phy_scan_tx2_out
PCIE_PHY_phy_scan_tx3_ana_dword_clk
PCIE_PHY_phy_scan_tx3_ana_dword_in
PCIE_PHY_phy_scan_tx3_ana_dword_out
PCIE_PHY_phy_scan_tx3_ana_word_clk
PCIE_PHY_phy_scan_tx3_ana_word_in
PCIE_PHY_phy_scan_tx3_ana_word_out
PCIE_PHY_phy_scan_tx3_in
PCIE_PHY_phy_scan_tx3_out
PCIE_PHY_phy_test_burnin
PCIE_PHY_phy_test_powerdown
PCIE_PHY_phy_test_stop_clk_en
PCIE_PHY_phy_tx0_flyover_data_m
PCIE_PHY_phy_tx0_flyover_data_p
PCIE_PHY_phy_tx1_flyover_data_m
PCIE_PHY_phy_tx1_flyover_data_p
PCIE_PHY_phy_tx2_flyover_data_m
PCIE_PHY_phy_tx2_flyover_data_p
PCIE_PHY_phy_tx3_flyover_data_m
PCIE_PHY_phy_tx3_flyover_data_p
PCIE_PHY_pipe_lane0_1_reset_n
PCIE_PHY_pipe_lane2_3_reset_n
PCIE_REF_DIG_CLK
PCIE_SUB_CON_x2_QACCEPTn_apb_aclk
PCIE_SUB_CON_x2_QACCEPTn_dbi_aclk
PCIE_SUB_CON_x2_QACCEPTn_mstr_aclk_slv_aclk
PCIE_SUB_CON_x2_QACTIVE_apb_aclk
PCIE_SUB_CON_x2_QACTIVE_dbi_aclk
PCIE_SUB_CON_x2_QACTIVE_mstr_aclk_slv_aclk
PCIE_SUB_CON_x2_QDENY_apb_aclk
PCIE_SUB_CON_x2_QDENY_dbi_aclk
PCIE_SUB_CON_x2_QDENY_mstr_aclk_slv_aclk
PCIE_SUB_CON_x2_QREQn_apb_aclk
PCIE_SUB_CON_x2_QREQn_dbi_aclk
PCIE_SUB_CON_x2_QREQn_mstr_aclk_slv_aclk
PCIE_SUB_CON_x2_TEST_AUXCLK
PCIE_SUB_CON_x2_TEST_MODE
PCIE_SUB_CON_x2_aux_clk_soc
PCIE_SUB_CON_x2_button_rst_n
PCIE_SUB_CON_x2_dbi_aclk_soc
PCIE_SUB_CON_x2_dbi_arready
PCIE_SUB_CON_x2_dbi_arvalid
PCIE_SUB_CON_x2_dbi_awready
PCIE_SUB_CON_x2_dbi_awvalid
PCIE_SUB_CON_x2_dbi_bready
PCIE_SUB_CON_x2_dbi_bvalid
PCIE_SUB_CON_x2_dbi_rlast
PCIE_SUB_CON_x2_dbi_rready
PCIE_SUB_CON_x2_dbi_rvalid
PCIE_SUB_CON_x2_dbi_wlast
PCIE_SUB_CON_x2_dbi_wready
PCIE_SUB_CON_x2_dbi_wvalid
PCIE_SUB_CON_x2_i_driver_apb_clk
PCIE_SUB_CON_x2_i_driver_apb_paddr
PCIE_SUB_CON_x2_i_driver_apb_penable
PCIE_SUB_CON_x2_i_driver_apb_psel
PCIE_SUB_CON_x2_i_driver_apb_pwdata
PCIE_SUB_CON_x2_i_driver_apb_pwrite
PCIE_SUB_CON_x2_i_driver_apb_rstn
PCIE_SUB_CON_x2_mstr_aclk_soc
PCIE_SUB_CON_x2_mstr_arready
PCIE_SUB_CON_x2_mstr_arvalid
PCIE_SUB_CON_x2_mstr_awready
PCIE_SUB_CON_x2_mstr_awvalid
PCIE_SUB_CON_x2_mstr_wready
PCIE_SUB_CON_x2_mstr_wvalid
PCIE_SUB_CON_x2_o_driver_apb_prdata
PCIE_SUB_CON_x2_o_driver_apb_pready
PCIE_SUB_CON_x2_o_driver_apb_pslverr
PCIE_SUB_CON_x2_pcie_irq
PCIE_SUB_CON_x2_perst_n
PCIE_SUB_CON_x2_phy_refclk_in
PCIE_SUB_CON_x2_power_up_rst_n
PCIE_SUB_CON_x2_slv_aclk_soc
PCIE_SUB_CON_x2_slv_arready
PCIE_SUB_CON_x2_slv_arvalid
PCIE_SUB_CON_x2_slv_awready
PCIE_SUB_CON_x2_slv_awvalid
PCIE_SUB_CON_x2_slv_bready
PCIE_SUB_CON_x2_slv_bvalid
PCIE_SUB_CON_x2_slv_rlast
PCIE_SUB_CON_x2_slv_rready
PCIE_SUB_CON_x2_slv_rvalid
PCIE_SUB_CON_x2_slv_wlast
PCIE_SUB_CON_x2_slv_wready
PCIE_SUB_CON_x2_slv_wvalid
PCIE_SUB_CON_x4_QACCEPTn_apb_aclk
PCIE_SUB_CON_x4_QACCEPTn_dbi_aclk
PCIE_SUB_CON_x4_QACCEPTn_mstr_aclk_slv_aclk
PCIE_SUB_CON_x4_QACTIVE_apb_aclk
PCIE_SUB_CON_x4_QACTIVE_dbi_aclk
PCIE_SUB_CON_x4_QACTIVE_mstr_aclk_slv_aclk
PCIE_SUB_CON_x4_QDENY_apb_aclk
PCIE_SUB_CON_x4_QDENY_dbi_aclk
PCIE_SUB_CON_x4_QDENY_mstr_aclk_slv_aclk
PCIE_SUB_CON_x4_QREQn_apb_aclk
PCIE_SUB_CON_x4_QREQn_dbi_aclk
PCIE_SUB_CON_x4_QREQn_mstr_aclk_slv_aclk
PCIE_SUB_CON_x4_TEST_AUXCLK
PCIE_SUB_CON_x4_TEST_MODE
PCIE_SUB_CON_x4_aux_clk_soc
PCIE_SUB_CON_x4_button_rst_n
PCIE_SUB_CON_x4_cr_para_sel
PCIE_SUB_CON_x4_dbi_aclk_soc
PCIE_SUB_CON_x4_dbi_arready
PCIE_SUB_CON_x4_dbi_arvalid
PCIE_SUB_CON_x4_dbi_awready
PCIE_SUB_CON_x4_dbi_awvalid
PCIE_SUB_CON_x4_dbi_bready
PCIE_SUB_CON_x4_dbi_bvalid
PCIE_SUB_CON_x4_dbi_rlast
PCIE_SUB_CON_x4_dbi_rready
PCIE_SUB_CON_x4_dbi_rvalid
PCIE_SUB_CON_x4_dbi_wlast
PCIE_SUB_CON_x4_dbi_wready
PCIE_SUB_CON_x4_dbi_wvalid
PCIE_SUB_CON_x4_ext_pclk_req
PCIE_SUB_CON_x4_i_driver_apb_clk
PCIE_SUB_CON_x4_i_driver_apb_paddr
PCIE_SUB_CON_x4_i_driver_apb_penable
PCIE_SUB_CON_x4_i_driver_apb_psel
PCIE_SUB_CON_x4_i_driver_apb_pwdata
PCIE_SUB_CON_x4_i_driver_apb_pwrite
PCIE_SUB_CON_x4_i_driver_apb_rstn
PCIE_SUB_CON_x4_mstr_aclk_soc
PCIE_SUB_CON_x4_mstr_arready
PCIE_SUB_CON_x4_mstr_arvalid
PCIE_SUB_CON_x4_mstr_awready
PCIE_SUB_CON_x4_mstr_awvalid
PCIE_SUB_CON_x4_mstr_wready
PCIE_SUB_CON_x4_mstr_wvalid
PCIE_SUB_CON_x4_o_driver_apb_prdata
PCIE_SUB_CON_x4_o_driver_apb_pready
PCIE_SUB_CON_x4_o_driver_apb_pslverr
PCIE_SUB_CON_x4_pcie_irq
PCIE_SUB_CON_x4_perst_n
PCIE_SUB_CON_x4_phy_lane0_rx2tx_par_lb_en
PCIE_SUB_CON_x4_phy_lane1_rx2tx_par_lb_en
PCIE_SUB_CON_x4_phy_lane2_rx2tx_par_lb_en
PCIE_SUB_CON_x4_phy_lane3_rx2tx_par_lb_en
PCIE_SUB_CON_x4_phy_refclk_in
PCIE_SUB_CON_x4_power_up_rst_n
PCIE_SUB_CON_x4_slv_aclk_soc
PCIE_SUB_CON_x4_slv_arready
PCIE_SUB_CON_x4_slv_arvalid
PCIE_SUB_CON_x4_slv_awready
PCIE_SUB_CON_x4_slv_awvalid
PCIE_SUB_CON_x4_slv_bready
PCIE_SUB_CON_x4_slv_bvalid
PCIE_SUB_CON_x4_slv_rlast
PCIE_SUB_CON_x4_slv_rready
PCIE_SUB_CON_x4_slv_rvalid
PCIE_SUB_CON_x4_slv_wlast
PCIE_SUB_CON_x4_slv_wready
PCIE_SUB_CON_x4_slv_wvalid
PCIE_SUB_CON_x4_sram_bypass
PIPE_MUX_PHY_MODE_SEL
