
// Connect ace_cluster_m
    assign ace_cluster_m.aclk             = /* FIXME */;
    assign ace_cluster_m.aresetn          = /* FIXME */;
    assign #100ps ace_cluster_m.acaddr           = AXI__ACADDR[43:0];
    assign #100ps ace_cluster_m.acprot           = AXI__ACPROT[2:0];
    assign #100ps ace_cluster_m.acsnoop          = AXI__ACSNOOP[3:0];
    assign #100ps ace_cluster_m.acvalid          = AXI__ACVALID;
    assign #100ps ace_cluster_m.arready          = AXI__ARREADY;
    assign #100ps ace_cluster_m.awready          = AXI__AWREADY;
    assign #100ps ace_cluster_m.bid              = AXI__BID[7:0];
    assign #100ps ace_cluster_m.bresp            = AXI__BRESP[1:0];
    assign #100ps ace_cluster_m.buser            = AXI__BUSER[0:0];
    assign #100ps ace_cluster_m.bvalid           = AXI__BVALID;
    assign #100ps ace_cluster_m.cdready          = AXI__CDREADY;
    assign #100ps ace_cluster_m.crready          = AXI__CRREADY;
    assign #100ps ace_cluster_m.rdata            = AXI__RDATA[127:0];
    assign #100ps ace_cluster_m.rid              = AXI__RID[8:0];
    assign #100ps ace_cluster_m.rlast            = AXI__RLAST;
    assign #100ps ace_cluster_m.rresp            = AXI__RRESP[3:0];
    assign #100ps ace_cluster_m.ruser            = AXI__RUSER[0:0];
    assign #100ps ace_cluster_m.rvalid           = AXI__RVALID;
    assign #100ps ace_cluster_m.wready           = AXI__WREADY;
    assign #100ps AXI__ACREADY                                       = ace_cluster_m.acready;
    assign #100ps AXI__ARADDR[43:0]                                  = ace_cluster_m.araddr;
    assign #100ps AXI__ARBAR[1:0]                                    = ace_cluster_m.arbar;
    assign #100ps AXI__ARBURST[1:0]                                  = ace_cluster_m.arburst;
    assign #100ps AXI__ARCACHE[3:0]                                  = ace_cluster_m.arcache;
    assign #100ps AXI__ARDOMAIN[1:0]                                 = ace_cluster_m.ardomain;
    assign #100ps AXI__ARID[8:0]                                     = ace_cluster_m.arid;
    assign #100ps AXI__ARLEN[7:0]                                    = ace_cluster_m.arlen;
    assign #100ps AXI__ARLOCK                                        = ace_cluster_m.arlock;
    assign #100ps AXI__ARPROT[2:0]                                   = ace_cluster_m.arprot;
    assign #100ps AXI__ARQOS[3:0]                                    = ace_cluster_m.arqos;
    assign #100ps AXI__ARREGION[3:0]                                 = ace_cluster_m.arregion;
    assign #100ps AXI__ARSIZE[2:0]                                   = ace_cluster_m.arsize;
    assign #100ps AXI__ARSNOOP[3:0]                                  = ace_cluster_m.arsnoop;
    assign #100ps AXI__ARUSER[7:0]                                   = ace_cluster_m.aruser;
    assign #100ps AXI__ARVALID                                       = ace_cluster_m.arvalid;
    assign #100ps AXI__AWADDR[43:0]                                  = ace_cluster_m.awaddr;
    assign #100ps AXI__AWBAR[1:0]                                    = ace_cluster_m.awbar;
    assign #100ps AXI__AWBURST[1:0]                                  = ace_cluster_m.awburst;
    assign #100ps AXI__AWCACHE[3:0]                                  = ace_cluster_m.awcache;
    assign #100ps AXI__AWDOMAIN[1:0]                                 = ace_cluster_m.awdomain;
    assign #100ps AXI__AWID[7:0]                                     = ace_cluster_m.awid;
    assign #100ps AXI__AWLEN[7:0]                                    = ace_cluster_m.awlen;
    assign #100ps AXI__AWLOCK                                        = ace_cluster_m.awlock;
    assign #100ps AXI__AWPROT[2:0]                                   = ace_cluster_m.awprot;
    assign #100ps AXI__AWQOS[3:0]                                    = ace_cluster_m.awqos;
    assign #100ps AXI__AWREGION[3:0]                                 = ace_cluster_m.awregion;
    assign #100ps AXI__AWSIZE[2:0]                                   = ace_cluster_m.awsize;
    assign #100ps AXI__AWSNOOP[2:0]                                  = ace_cluster_m.awsnoop;
    assign #100ps /* FIXME */                                        = ace_cluster_m.awunique;
    assign #100ps AXI__AWUSER[7:0]                                   = ace_cluster_m.awuser;
    assign #100ps AXI__AWVALID                                       = ace_cluster_m.awvalid;
    assign #100ps AXI__BREADY                                        = ace_cluster_m.bready;
    assign #100ps AXI__CDDATA[127:0]                                 = ace_cluster_m.cddata;
    assign #100ps AXI__CDLAST                                        = ace_cluster_m.cdlast;
    assign #100ps AXI__CDVALID                                       = ace_cluster_m.cdvalid;
    assign #100ps AXI__CRRESP[4:0]                                   = ace_cluster_m.crresp;
    assign #100ps AXI__CRVALID                                       = ace_cluster_m.crvalid;
    assign #100ps AXI__RACK                                          = ace_cluster_m.rack;
    assign #100ps AXI__RREADY                                        = ace_cluster_m.rready;
    assign #100ps AXI__WACK                                          = ace_cluster_m.wack;
    assign #100ps AXI__WDATA[127:0]                                  = ace_cluster_m.wdata;
    assign #100ps AXI__WLAST                                         = ace_cluster_m.wlast;
    assign #100ps AXI__WSTRB[15:0]                                   = ace_cluster_m.wstrb;
    assign #100ps AXI__WUSER[0:0]                                    = ace_cluster_m.wuser;
    assign #100ps AXI__WVALID                                        = ace_cluster_m.wvalid;
